library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity memory is
Port ( 
	dir : in STD_LOGIC_VECTOR (11 downto 0);
	data : out STD_LOGIC_VECTOR (93 downto 0));
end memory;

architecture Behavioral of memory is

begin
	process(dir)
	begin
	
		-- DATA FORMAT
		-- |    PRUEBA    |VF| Ins |                LIGA                 |
		--  P4 P3 P2 P1 P0 VF I1 I0 L11 L10 L9 L8 L7 L6 L5 L4 L3 L2 L1 L0 nCRI EB1 EB0 nWB EA1 EA0 nWA selbus UPA9 UPA8 UPA7 UPA6 UPA5 UPA4 UPA3 UPA2 UPA1 UPA0 nOEUPA nDUPA selmux nEX2 nEX1 nEX0 X2 X1 X0 EnaY nERA2 nERA1 nERA0 RA2 RA1 RA0 nEAP2 nEAP1 nEAP0 AP2 AP1 AP0 nEPC2 nEPC1 nEPC0 PC2 PC1 PC0 nCBD nAS nRW BD DINT HINT SET_IRQ SET_XIRQ B9 B8 B7 B6 B5 B4 B3 B2 B1 B0 CC CN CV CZ CI CH CX CS nHB ACCSEC

		-- Cadena por default: "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010"
		
		--if(dir=    X"000") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010";
		--elsif(dir= X"001") then data <= "00000" & "0" & "00" & "000000000000" & "00000000000000000000000000000000000000000000000000000000000000000000000000"; 
												  
												  
		if(dir=    X"000") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"001") then data <= "00000" & "0" & "00" & "000000000000" & "00010010000000000011011100001110001110001110011010000000000000000000000010";
		elsif(dir= X"002") then data <= "00000" & "0" & "10" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010";		
		
		elsif(dir= X"860") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"861") then data <= "00000" & "0" & "00" & "000000000000" & "10010100000000000011011100001110001110001110011010000000000000000000000010";
		elsif(dir= X"862") then data <= "01111" & "1" & "11" & "000000000000" & "10010010000000000011011100001110001110001110001110000000010011000111000010";
		elsif(dir= X"863") then data <= "11000" & "0" & "01" & "000000000001" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		
		elsif(dir= X"C60") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"C61") then data <= "00000" & "0" & "00" & "000000000000" & "10100010000000000011011100001110001110001110011010000000000000000000000010";
		elsif(dir= X"C62") then data <= "01111" & "1" & "11" & "000000000000" & "10010010000000000011011100001110001110001110001110000000100101000111000010";
		elsif(dir= X"C63") then data <= "11000" & "0" & "01" & "000000000001" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		
		elsif(dir= X"180") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100011110001110000110000110000000000000000000000010";
		elsif(dir= X"181") then data <= "00000" & "0" & "00" & "000000000000" & "00010010000000000011011100001110001110001110011010000000000000000000000010";
		elsif(dir= X"182") then data <= "00000" & "0" & "10" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010";
		
		elsif(dir= X"CE0") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"CE1") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011010110001110001110001110011011000000000000000000000010";
		elsif(dir= X"CE2") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"CE3") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011001101110001110001110011010000000000000000000000010";
		elsif(dir= X"CE4") then data <= "01111" & "1" & "11" & "000000000000" & "10010010000000000011011100001110001110001110001110000000110111000111000010";
		elsif(dir= X"CE5") then data <= "11000" & "0" & "01" & "000000000001" & "10010010000000000011011100001110001110000110000110000000000000000000000010";

	
		
		elsif(dir= X"1B0") then data <= "00000" & "0" & "00" & "000000000000" & "11111110000000000111111100001110001110001110001110000000000000000000000010";
		elsif(dir= X"1B1") then data <= "01111" & "1" & "11" & "000000000000" & "10010100000000000000011100001110001110001110001110000000000000001111010010";
		elsif(dir= X"1B2") then data <= "11000" & "0" & "01" & "000000000001" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
	
		elsif(dir= X"7E0") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"7E1") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001011001110001110011011000000000000000000000010";
		elsif(dir= X"7E2") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"7E3") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001100111110001110011010000000000000000000000010";
		elsif(dir= X"7E4") then data <= "01111" & "1" & "11" & "000000000000" & "10010010000000000011011100001000001110001001011110000000000000000000000010";
		elsif(dir= X"7E5") then data <= "11000" & "0" & "01" & "000000000001" & "10010010000000000011011100001110001110000110000110000000000000000000000010";
		else data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010"; -- Default
		end if;
	end process;
end Behavioral;